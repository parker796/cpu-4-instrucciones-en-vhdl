library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity lcd is
    port(
        clk_50:in std_logic;
        numins:in std_logic_vector(3 downto 0);
        palabra:out std_logic_vector(12 downto 0)
    );
end entity lcd;

architecture beh of lcd is
    signal clk:std_logic:= '0';
    signal comandos:natural range 0 to 5;
    signal load1:natural range 0 to 27;
    signal load2:natural range 0 to 23;
    signal add:natural range 0 to 31;
    signal mov:natural range 0 to 27;
    signal sub:natural range 0 to 31;
    --en esta parte hacemos la deteccion de un flanco para controlar el tiempo que en este caso son 100000 milisegundo
begin
    process(clk_50)
        variable cuenta:natural range 0 to 100_000 :=0 ;
    begin   
        if clk_50'event and clk_50 = '1' then
            cuenta := cuenta + 1;
            if cuenta = 100_000 then 
                cuenta := 0;
                clk <= not clk;
            end if;
        end if;
    end process;

    process(clk)
    begin
        if clk'event and clk = '1' then
            case comandos is
                when 0 =>
                    palabra <= "1110000000001";
                    comandos  <= comandos + 1;
                when 1 =>
                    palabra <= "1100000000110";
                    comandos  <= comandos + 1;
                when 2 =>
                    palabra <= "1110000001111";
                    comandos  <= comandos + 1;
                when 3 =>
                    palabra <= "1100001110000";
                    comandos  <= comandos + 1;
                when 4 => 
                    palabra <= "1110000111000";
                    comandos  <= comandos + 1;

                when 5 =>
                    case numins is
                        when "0000" =>
                            case load1 is
                                when 0 =>
                                    palabra <= "1101001101100";
                                    load1  <= load1 + 1;
                                when 1 =>
                                    palabra <= "1111001101100";
                                    load1  <= load1 + 1;
                                when 2 =>
                                    palabra <= "1101001101111";
                                    load1  <= load1 + 1;
                                when 3 =>
                                    palabra <= "1111001101111";
                                    load1  <= load1 + 1;
                                when 4 =>
                                    palabra <= "1101001100001";
                                    load1  <= load1 + 1;
                                when 5 =>
                                    palabra <= "1111001100001";
                                    load1  <= load1 + 1;
                                when 6 =>
                                    palabra <= "1101001100100";
                                    load1  <= load1 + 1;
                                when 7 =>
                                    palabra <= "1111001100100";
                                    load1  <= load1 + 1;
                                when 8 =>
                                    palabra <= "1101000100000";
                                    load1  <= load1 + 1;
                                when 9 =>
                                    palabra <= "1111000100000";
                                    load1  <= load1 + 1;
                                when 10 =>
                                    palabra <= "1101000110000";
                                    load1  <= load1 + 1;
                                when 11 =>
                                    palabra <= "1111000110000";
                                    load1  <= load1 + 1;
                                when 12 =>
                                    palabra <= "1101001111000";
                                    load1  <= load1 + 1;
                                when 13 =>
                                    palabra <= "1111001111000";
                                    load1  <= load1 + 1;
                                when 14 =>
                                    palabra <= "1101001000001";
                                    load1  <= load1 + 1;
                                when 15 =>
                                    palabra <= "1111001000001";
                                    load1  <= load1 + 1;
                                when 16 =>
                                    palabra <= "1101000101100";
                                    load1  <= load1 + 1;
                                when 17 =>
                                    palabra <= "1111000101100";
                                    load1  <= load1 + 1;
                                when 18 =>
                                    palabra <= "1101000100000";
                                    load1  <= load1 + 1;
                                when 19 =>
                                    palabra <= "1111000100000";
                                    load1  <= load1 + 1;
                                when 20 =>
                                    palabra <= "1101000100101";
                                    load1  <= load1 + 1;
                                when 21 =>
                                    palabra <= "1111000100101";
                                    load1  <= load1 + 1;
                                when 22 =>
                                    palabra <= "1101001110010";
                                    load1  <= load1 + 1;
                                when 23 =>
                                    palabra <= "1111001110010";
                                    load1  <= load1 + 1;
                                when 24 =>
                                    palabra <= "1101000110000";
                                    load1  <= load1 + 1;
                                when 25 =>
                                    palabra <= "1111000110000";
                                    load1  <= load1 + 1;
                                when 26 =>
                                    palabra <= "1101000100000";
                                    load1  <= load1 + 1;
                                when 27 =>
                                    palabra <= "1110000000001";
                            end case;
                        when "0001" =>
                            case load2 is
                                when 0 =>
                                    palabra <= "1101001101100";
                                    load2  <= load2 + 1;
                                when 1 =>
                                    palabra <= "1111001101100";
                                    load2  <= load2 + 1;
                                when 2 =>
                                    palabra <= "1101001101111";
                                    load2  <= load2 + 1;
                                when 3 =>
                                    palabra <= "1111001101111";
                                    load2  <= load2 + 1;
                                when 4 =>
                                    palabra <= "1101001100001";
                                    load2  <= load2 + 1;
                                when 5 =>
                                    palabra <= "1111001100001";
                                    load2  <= load2 + 1;
                                when 6 =>
                                    palabra <= "1101001100100";
                                    load2  <= load2 + 1;
                                when 7 =>
                                    palabra <= "1111001100100";
                                    load2  <= load2 + 1;
                                when 8 =>
                                    palabra <= "1101000100000";
                                    load2  <= load2 + 1;
                                when 9 =>
                                    palabra <= "1111000100000";
                                    load2  <= load2 + 1;
                                when 10 =>
                                    palabra <= "1101000110011";
                                    load2  <= load2 + 1;
                                when 11 =>
                                    palabra <= "1111000110011";
                                    load2  <= load2 + 1;
                                when 12 =>
                                    palabra <= "1101000101100";
                                    load2  <= load2 + 1;
                                when 13 =>
                                    palabra <= "1111000101100";
                                    load2  <= load2 + 1;
                                when 14 =>
                                    palabra <= "1101000100000";
                                    load2  <= load2 + 1;
                                when 15 =>
                                    palabra <= "1111000100000";
                                    load2  <= load2 + 1;
                                when 16 =>
                                    palabra <= "1101000100101";
                                    load2  <= load2 + 1;
                                when 17 =>
                                    palabra <= "1111000100101";
                                    load2  <= load2 + 1;
                                when 18 =>
                                    palabra <= "1101001110010";
                                    load2  <= load2 + 1;
                                when 19 =>
                                    palabra <= "1111001110010";
                                    load2  <= load2 + 1;
                                when 20 =>
                                    palabra <= "1101000110001";
                                    load2  <= load2 + 1;
                                when 21 =>
                                    palabra <= "1111000110001";
                                    load2  <= load2 + 1;
                                when 22 =>
                                    palabra <= "1101000100000";
                                    load2  <= load2 + 1;
                                when 23 =>
                                    palabra <= "1110000000001"; 
                            end case;
                        when "0010" =>
                            case add is
                                when 0 =>
                                    palabra <= "1101001100001";
                                    add  <= add + 1;
                                when 1 =>
                                    palabra <= "1111001100001";
                                    add  <= add + 1;
                                when 2 =>
                                    palabra <= "1101001100100";
                                    add  <= add + 1;
                                when 3 =>
                                    palabra <= "1111001100100";
                                    add  <= add + 1;
                                when 4 =>
                                    palabra <= "1101001100100";
                                    add  <= add + 1;
                                when 5 =>
                                    palabra <= "1111001100100";
                                    add  <= add + 1;
                                when 6 =>
                                    palabra <= "1101000100000";
                                    add  <= add + 1;
                                when 7 =>
                                    palabra <= "1111000100000";
                                    add  <= add + 1;
                                when 8 =>
                                    palabra <= "1101000100101";
                                    add  <= add + 1;
                                when 9 =>
                                    palabra <= "1111000100101";
                                    add  <= add + 1;
                                when 10 =>
                                    palabra <= "1101001110010";
                                    add  <= add + 1;
                                when 11 =>
                                    palabra <= "1111001110010";
                                    add  <= add + 1;
                                when 12 =>
                                    palabra <= "1101000110000";
                                    add  <= add + 1;
                                when 13 =>
                                    palabra <= "1111000110000";
                                    add  <= add + 1;
                                when 14 =>
                                    palabra <= "1101000101100";
                                    add  <= add + 1;
                                when 15 =>
                                    palabra <= "1111000101100";
                                    add  <= add + 1;
                                when 16 =>
                                    palabra <= "1101000100101";
                                    add  <= add + 1;
                                when 17 =>
                                    palabra <= "1111000100101";
                                    add  <= add + 1;
                                when 18 =>
                                    palabra <= "1101001110010";
                                    add  <= add + 1;
                                when 19 =>
                                    palabra <= "1111001110010";
                                    add  <= add + 1;
                                when 20 =>
                                    palabra <= "1101000110001";
                                    add  <= add + 1;
                                when 21 =>
                                    palabra <= "1111000110001"; 
                                    add  <= add + 1;
                                when 22 =>
                                    palabra <= "1101000101100";
                                    add  <= add + 1;
                                when 23 =>
                                    palabra <= "1111000101100";
                                    add  <= add + 1;
                                when 24 =>
                                    palabra <= "1101000100101";
                                    add  <= add + 1;
                                when 25 =>
                                    palabra <= "1111000100101";
                                    add  <= add + 1;
                                when 26 =>
                                    palabra <= "1101001110010";
                                    add  <= add + 1;
                                when 27 =>
                                    palabra <= "1111001110010";
                                    add  <= add + 1;
                                when 28 =>
                                    palabra <= "1101000110010";
                                    add  <= add + 1;
                                when 29 =>
                                    palabra <= "1111000110010"; 
                                    add  <= add + 1;
                                when 30 =>
                                    palabra <= "1101000110010";
                                    add  <= add + 1;
                                when 31 =>
                                    palabra <= "1110000000001"; 
                            end case;
                        when "0011" =>
                            case mov is
                            when 0 =>
                                palabra <= "1101001101101";
                                mov  <= mov + 1;
                            when 1 =>
                                palabra <= "1111001101101";
                                mov  <= mov + 1;
                            when 2 =>
                                palabra <= "1101001101111";
                                mov  <= mov + 1;
                            when 3 =>
                                palabra <= "1111001101111";
                                mov  <= mov + 1;
                            when 4 =>
                                palabra <= "1101001110110";
                                mov  <= mov + 1;
                            when 5 =>
                                palabra <= "1111001110110";
                                mov  <= mov + 1;
                            when 6 =>
                                palabra <= "1101001100101";
                                mov  <= mov + 1;
                            when 7 =>
                                palabra <= "1111001100101";
                                mov  <= mov + 1;
                            when 8 =>
                                palabra <= "1101000100000";
                                mov  <= mov + 1;
                            when 9 =>
                                palabra <= "1111000100000";
                                mov  <= mov + 1;
                            when 10 =>
                                palabra <= "1101000100101";
                                mov  <= mov + 1;
                            when 11 =>
                                palabra <= "1111000100101";
                                mov  <= mov + 1;
                            when 12 =>
                                palabra <= "1101001110010";
                                mov  <= mov + 1;
                            when 13 =>
                                palabra <= "1111001110010";
                                mov  <= mov + 1;
                            when 14 =>
                                palabra <= "1101000110010";
                                mov  <= mov + 1;
                            when 15 =>
                                palabra <= "1111000110010";
                                mov  <= mov + 1;
                            when 16 =>
                                palabra <= "1101000101100";
                                mov  <= mov + 1;
                            when 17 =>
                                palabra <= "1111000101100";
                                mov  <= mov + 1;
                            when 18 =>
                                palabra <= "1101000100000";
                                mov  <= mov + 1;
                            when 19 =>
                                palabra <= "1111000100000";
                                mov  <= mov + 1;
                            when 20 =>
                                palabra <= "1101000100101";
                                mov  <= mov + 1;
                            when 21 =>
                                palabra <= "1111000100101"; 
                                mov  <= mov + 1;
                            when 22 =>
                                palabra <= "1101001110010";
                                mov  <= mov + 1;
                            when 23 =>
                                palabra <= "1111001110010";
                                mov  <= mov + 1;
                            when 24 =>
                                palabra <= "1101000110011";
                                mov  <= mov + 1;
                            when 25 =>
                                palabra <= "1111000110011";
                                mov  <= mov + 1;
                            when 26 =>
                                palabra <= "1101000100000";
                                mov  <= mov + 1;
                            when 27 =>
                                palabra <= "1110000000001";
                        end case;
                    when "0100" =>
                        case sub is
                        when 0 =>
                            palabra <= "1101001110011";
                            sub  <= sub + 1;
                        when 1 =>
                            palabra <= "1111001110011";
                            sub  <= sub + 1;
                        when 2 =>
                            palabra <= "1101001110101";
                            sub  <= sub + 1;
                        when 3 =>
                            palabra <= "1111001110101";
                            sub  <= sub + 1;
                        when 4 =>
                            palabra <= "1101001100010";
                            sub  <= sub + 1;
                        when 5 =>
                            palabra <= "1111001100010";
                            sub  <= sub + 1;
                        when 6 =>
                            palabra <= "1101000100000";
                            sub  <= sub + 1;
                        when 7 =>
                            palabra <= "1111000100000";
                            sub  <= sub + 1;
                        when 8 =>
                            palabra <= "1101000100101";
                            sub  <= sub + 1;
                        when 9 =>
                            palabra <= "1111000100101";
                            sub  <= sub + 1;
                        when 10 =>
                            palabra <= "1101001110010";
                            sub  <= sub + 1;
                        when 11 =>
                            palabra <= "1111001110010";
                            sub  <= sub + 1;
                        when 12 =>
                            palabra <= "1101000110011";
                            sub  <= sub + 1;
                        when 13 =>
                            palabra <= "1111000110011";
                            sub  <= sub + 1;
                        when 14 =>
                            palabra <= "1101000101100";
                            sub  <= sub + 1;
                        when 15 =>
                            palabra <= "1111000101100";
                            sub  <= sub + 1;
                        when 16 =>
                            palabra <= "1101000100101";
                            sub  <= sub + 1;
                        when 17 =>
                            palabra <= "1111000100101";
                            sub  <= sub + 1;
                        when 18 =>
                            palabra <= "1101001110010";
                            sub  <= sub + 1;
                        when 19 =>
                            palabra <= "1111001110010";
                            sub  <= sub + 1;
                        when 20 =>
                            palabra <= "1101000110000";
                            sub  <= sub + 1;
                        when 21 =>
                            palabra <= "1111000110000"; 
                            sub  <= sub + 1;
                        when 22 =>
                            palabra <= "1101000101100";
                            sub  <= sub + 1;
                        when 23 =>
                            palabra <= "1111000101100";
                            sub  <= sub + 1;
                        when 24 =>
                            palabra <= "1101000100101";
                            sub  <= sub + 1;
                        when 25 =>
                            palabra <= "1111000100101";
                            sub  <= sub + 1;
                        when 26 =>
                            palabra <= "1101001110010";
                            sub  <= sub + 1;
                        when 27 =>
                            palabra <= "1111001110010";
                            sub  <= sub + 1;
                        when 28 =>
                            palabra <= "1101000110001";
                            sub  <= sub + 1;
                        when 29 =>
                            palabra <= "1111000110001"; 
                            sub  <= sub + 1;
                        when 30 =>
                            palabra <= "1101000110010";
                            sub  <= sub + 1;
                        when 31 =>
                            palabra <= "1110000000001";
                        end case;
                    when others =>
                    end case;
                end case;
        end if;
    end process;
end architecture beh;
